module ROM #(
    MemSize = 1024
) (
    input                   clk_i,
    input                   ctrlSignal_i,
    input       [31:0]      addrwire_i, // ��д��ַ
    output  reg [31:0]      data_o
);

reg [7:0]   mm[MemSize - 1 : 0];

integer n;
initial begin
	{ mm[ 3], mm[ 2], mm[ 1], mm[ 0] } = 32'b000000000001_00000_000_00011_0010011;
	{ mm[ 7], mm[ 6], mm[ 5], mm[ 4] } = 32'b000000000001_00000_000_00100_0010011;
	{ mm[11], mm[10], mm[ 9], mm[ 8] } = 32'b000000000010_00000_000_00101_0010011;
	{ mm[15], mm[14], mm[13], mm[12] } = 32'b000000110010_00000_000_00110_0010011;
	{ mm[19], mm[18], mm[17], mm[16] } = 32'b111111111101_00110_000_00110_0010011;
	{ mm[23], mm[22], mm[21], mm[20] } = 32'b000000000000_00100_000_00011_0010011;
	{ mm[27], mm[26], mm[25], mm[24] } = 32'b000000000000_00101_000_00100_0010011;
	{ mm[31], mm[30], mm[29], mm[28] } = 32'b0000000_00100_00011_000_00101_0110011;
	{ mm[35], mm[34], mm[33], mm[32] } = 32'b111111111111_00110_000_00110_0010011;
	{ mm[39], mm[38], mm[37], mm[36] } = 32'b1111111_00110_00000_100_10001_1100011;
	{ mm[43], mm[42], mm[41], mm[40] } = 32'b0000000_00101_00000_100_00100_0100011;
	{ mm[47], mm[46], mm[45], mm[44] } = 32'b000000000100_00000_100_00111_0000011;
	{ mm[51], mm[50], mm[49], mm[48] } = 32'b00000000100000000000_00100_1101111;
	{ mm[55], mm[54], mm[53], mm[52] } = 32'b1111111_00000_00000_000_11101_1100011;
	{ mm[59], mm[58], mm[57], mm[56] } = 32'b000000000000_00100_000_00000_1100111;

    for (n = 60; n < MemSize; n = n + 1) begin
        mm[n] <= {8{1'b0}};
    end
end

wire    [31:0]  addr0;
wire    [31:0]  addr1;
wire    [31:0]  addr2;
wire    [31:0]  addr3;

assign  addr0   =   { addrwire_i[31:2], 2'b00 };
assign  addr1   =   { addrwire_i[31:2], 2'b01 };
assign  addr2   =   { addrwire_i[31:2], 2'b10 };
assign  addr3   =   { addrwire_i[31:2], 2'b11 };

always @(posedge clk_i) begin
    if (ctrlSignal_i)
        data_o  <=  { mm[addr3],  mm[addr2], mm[addr1],  mm[addr0] };
    else 
        data_o  <=  32'b0;
end   

endmodule